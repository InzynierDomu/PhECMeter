.title KiCad schematic
A1 NC_01 NC_02 NC_03 GND Net-_A1-Pad5_ Net-_A1-Pad6_ NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 Arduino_Nano_v3.x
SW1 GND Net-_A1-Pad5_ SW_Push
SW2 GND Net-_A1-Pad6_ SW_Push
.end
